// SPDX-FileCopyrightText: 2022 CERN (home.cern)
//
// SPDX-License-Identifier: CERN-OHL-W-2.0+

`define ADDR_FD_DCR                    6'h0
`define FD_DCR_ENABLE_OFFSET 0
`define FD_DCR_ENABLE 32'h00000001
`define FD_DCR_MODE_OFFSET 1
`define FD_DCR_MODE 32'h00000002
`define FD_DCR_PG_ARM_OFFSET 2
`define FD_DCR_PG_ARM 32'h00000004
`define FD_DCR_PG_TRIG_OFFSET 3
`define FD_DCR_PG_TRIG 32'h00000008
`define FD_DCR_UPDATE_OFFSET 4
`define FD_DCR_UPDATE 32'h00000010
`define FD_DCR_UPD_DONE_OFFSET 5
`define FD_DCR_UPD_DONE 32'h00000020
`define FD_DCR_FORCE_DLY_OFFSET 6
`define FD_DCR_FORCE_DLY 32'h00000040
`define FD_DCR_NO_FINE_OFFSET 7
`define FD_DCR_NO_FINE 32'h00000080
`define FD_DCR_FORCE_HI_OFFSET 8
`define FD_DCR_FORCE_HI 32'h00000100
`define ADDR_FD_FRR                    6'h4
`define ADDR_FD_U_STARTH               6'h8
`define ADDR_FD_U_STARTL               6'hc
`define ADDR_FD_C_START                6'h10
`define ADDR_FD_F_START                6'h14
`define ADDR_FD_U_ENDH                 6'h18
`define ADDR_FD_U_ENDL                 6'h1c
`define ADDR_FD_C_END                  6'h20
`define ADDR_FD_F_END                  6'h24
`define ADDR_FD_U_DELTA                6'h28
`define ADDR_FD_C_DELTA                6'h2c
`define ADDR_FD_F_DELTA                6'h30
`define ADDR_FD_RCR                    6'h34
`define FD_RCR_REP_CNT_OFFSET 0
`define FD_RCR_REP_CNT 32'h0000ffff
`define FD_RCR_CONT_OFFSET 16
`define FD_RCR_CONT 32'h00010000
