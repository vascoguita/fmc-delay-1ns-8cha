-- SPDX-FileCopyrightText: 2022 CERN (home.cern)
--
-- SPDX-License-Identifier: CERN-OHL-W-2.0+

---------------------------------------------------------------------------------------
-- Title          : Wishbone slave core for Fine Delay Channel WB Slave
---------------------------------------------------------------------------------------
-- File           : fd_channel_wbgen2_pkg.vhd
-- Author         : auto-generated by wbgen2 from fd_channel_wishbone_slave.wb
-- Created        : Wed Mar 20 23:27:12 2019
-- Standard       : VHDL'87
---------------------------------------------------------------------------------------
-- THIS FILE WAS GENERATED BY wbgen2 FROM SOURCE FILE fd_channel_wishbone_slave.wb
-- DO NOT HAND-EDIT UNLESS IT'S ABSOLUTELY NECESSARY!
---------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package fd_channel_wbgen2_pkg is
  
  
  -- Input registers (user design -> WB slave)
  
  type t_fd_channel_in_registers is record
    dcr_pg_trig_i                            : std_logic;
    dcr_upd_done_i                           : std_logic;
  end record;
  
  constant c_fd_channel_in_registers_init_value: t_fd_channel_in_registers := (
    dcr_pg_trig_i => '0',
    dcr_upd_done_i => '0'
  );
  
  -- Output registers (WB slave -> user design)
  
  type t_fd_channel_out_registers is record
    dcr_enable_o                             : std_logic;
    dcr_mode_o                               : std_logic;
    dcr_pg_arm_o                             : std_logic;
    dcr_update_o                             : std_logic;
    dcr_force_dly_o                          : std_logic;
    dcr_no_fine_o                            : std_logic;
    dcr_force_hi_o                           : std_logic;
    frr_o                                    : std_logic_vector(9 downto 0);
    u_starth_o                               : std_logic_vector(7 downto 0);
    u_startl_o                               : std_logic_vector(31 downto 0);
    c_start_o                                : std_logic_vector(27 downto 0);
    f_start_o                                : std_logic_vector(11 downto 0);
    u_endh_o                                 : std_logic_vector(7 downto 0);
    u_endl_o                                 : std_logic_vector(31 downto 0);
    c_end_o                                  : std_logic_vector(27 downto 0);
    f_end_o                                  : std_logic_vector(11 downto 0);
    u_delta_o                                : std_logic_vector(3 downto 0);
    c_delta_o                                : std_logic_vector(27 downto 0);
    f_delta_o                                : std_logic_vector(11 downto 0);
    rcr_rep_cnt_o                            : std_logic_vector(15 downto 0);
    rcr_cont_o                               : std_logic;
  end record;
  
  constant c_fd_channel_out_registers_init_value: t_fd_channel_out_registers := (
    dcr_enable_o => '0',
    dcr_mode_o => '0',
    dcr_pg_arm_o => '0',
    dcr_update_o => '0',
    dcr_force_dly_o => '0',
    dcr_no_fine_o => '0',
    dcr_force_hi_o => '0',
    frr_o => (others => '0'),
    u_starth_o => (others => '0'),
    u_startl_o => (others => '0'),
    c_start_o => (others => '0'),
    f_start_o => (others => '0'),
    u_endh_o => (others => '0'),
    u_endl_o => (others => '0'),
    c_end_o => (others => '0'),
    f_end_o => (others => '0'),
    u_delta_o => (others => '0'),
    c_delta_o => (others => '0'),
    f_delta_o => (others => '0'),
    rcr_rep_cnt_o => (others => '0'),
    rcr_cont_o => '0'
  );

function "or" (left, right: t_fd_channel_in_registers) return t_fd_channel_in_registers;
function f_x_to_zero (x:std_logic) return std_logic;
function f_x_to_zero (x:std_logic_vector) return std_logic_vector;

component fd_channel_wb_slave is
  port (
    rst_n_i                                  : in     std_logic;
    clk_sys_i                                : in     std_logic;
    wb_adr_i                                 : in     std_logic_vector(3 downto 0);
    wb_dat_i                                 : in     std_logic_vector(31 downto 0);
    wb_dat_o                                 : out    std_logic_vector(31 downto 0);
    wb_cyc_i                                 : in     std_logic;
    wb_sel_i                                 : in     std_logic_vector(3 downto 0);
    wb_stb_i                                 : in     std_logic;
    wb_we_i                                  : in     std_logic;
    wb_ack_o                                 : out    std_logic;
    wb_err_o                                 : out    std_logic;
    wb_rty_o                                 : out    std_logic;
    wb_stall_o                               : out    std_logic;
    clk_ref_i                                : in     std_logic;
    regs_i                                   : in     t_fd_channel_in_registers;
    regs_o                                   : out    t_fd_channel_out_registers
  );
end component;

end package;

package body fd_channel_wbgen2_pkg is
function f_x_to_zero (x:std_logic) return std_logic is
begin
  if x = '1' then
    return '1';
  else
    return '0';
  end if;
end function;

function f_x_to_zero (x:std_logic_vector) return std_logic_vector is
  variable tmp: std_logic_vector(x'length-1 downto 0);
begin
  for i in 0 to x'length-1 loop
    if(x(i) = 'X' or x(i) = 'U') then
      tmp(i):= '0';
    else
      tmp(i):=x(i);
    end if; 
  end loop; 
  return tmp;
end function;

function "or" (left, right: t_fd_channel_in_registers) return t_fd_channel_in_registers is
  variable tmp: t_fd_channel_in_registers;
begin
  tmp.dcr_pg_trig_i := f_x_to_zero(left.dcr_pg_trig_i) or f_x_to_zero(right.dcr_pg_trig_i);
  tmp.dcr_upd_done_i := f_x_to_zero(left.dcr_upd_done_i) or f_x_to_zero(right.dcr_upd_done_i);
  return tmp;
end function;

end package body;
