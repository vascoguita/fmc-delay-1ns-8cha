-- SPDX-FileCopyrightText: 2022 CERN (home.cern)
--
-- SPDX-License-Identifier: CERN-OHL-W-2.0+

---------------------------------------------------------------------------------------
-- Title          : Wishbone slave core for Fine Delay Main WB Slave
---------------------------------------------------------------------------------------
-- File           : fd_main_wishbone_slave.vhd
-- Author         : auto-generated by wbgen2 from fd_main_wishbone_slave.wb
-- Created        : Thu May 28 16:19:19 2020
-- Standard       : VHDL'87
---------------------------------------------------------------------------------------
-- THIS FILE WAS GENERATED BY wbgen2 FROM SOURCE FILE fd_main_wishbone_slave.wb
-- DO NOT HAND-EDIT UNLESS IT'S ABSOLUTELY NECESSARY!
---------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.wbgen2_pkg.all;

use work.fd_main_wbgen2_pkg.all;


entity fd_main_wb_slave is
port (
  rst_n_i                                  : in     std_logic;
  clk_sys_i                                : in     std_logic;
  wb_adr_i                                 : in     std_logic_vector(5 downto 0);
  wb_dat_i                                 : in     std_logic_vector(31 downto 0);
  wb_dat_o                                 : out    std_logic_vector(31 downto 0);
  wb_cyc_i                                 : in     std_logic;
  wb_sel_i                                 : in     std_logic_vector(3 downto 0);
  wb_stb_i                                 : in     std_logic;
  wb_we_i                                  : in     std_logic;
  wb_ack_o                                 : out    std_logic;
  wb_err_o                                 : out    std_logic;
  wb_rty_o                                 : out    std_logic;
  wb_stall_o                               : out    std_logic;
  wb_int_o                                 : out    std_logic;
  clk_ref_i                                : in     std_logic;
  tcr_rd_ack_o                             : out    std_logic;
  dmtr_in_rd_ack_o                         : out    std_logic;
  dmtr_out_rd_ack_o                        : out    std_logic;
  tsbcr_read_ack_o                         : out    std_logic;
  fid_read_ack_o                           : out    std_logic;
  irq_ts_buf_notempty_i                    : in     std_logic;
  irq_dmtd_spll_i                          : in     std_logic;
  irq_sync_status_i                        : in     std_logic;
  regs_i                                   : in     t_fd_main_in_registers;
  regs_o                                   : out    t_fd_main_out_registers
);
end fd_main_wb_slave;

architecture syn of fd_main_wb_slave is

signal fd_main_gcr_bypass_int                   : std_logic      ;
signal fd_main_gcr_bypass_sync0                 : std_logic      ;
signal fd_main_gcr_bypass_sync1                 : std_logic      ;
signal fd_main_gcr_input_en_int                 : std_logic      ;
signal fd_main_gcr_input_en_sync0               : std_logic      ;
signal fd_main_gcr_input_en_sync1               : std_logic      ;
signal fd_main_tcr_wr_enable_int                : std_logic      ;
signal fd_main_tcr_cap_time_int                 : std_logic      ;
signal fd_main_tcr_cap_time_int_delay           : std_logic      ;
signal fd_main_tcr_cap_time_sync0               : std_logic      ;
signal fd_main_tcr_cap_time_sync1               : std_logic      ;
signal fd_main_tcr_cap_time_sync2               : std_logic      ;
signal fd_main_tcr_set_time_int                 : std_logic      ;
signal fd_main_tcr_set_time_int_delay           : std_logic      ;
signal fd_main_tcr_set_time_sync0               : std_logic      ;
signal fd_main_tcr_set_time_sync1               : std_logic      ;
signal fd_main_tcr_set_time_sync2               : std_logic      ;
signal fd_main_tm_sech_int_read                 : std_logic_vector(7 downto 0);
signal fd_main_tm_sech_int_write                : std_logic_vector(7 downto 0);
signal fd_main_tm_sech_lw                       : std_logic      ;
signal fd_main_tm_sech_lw_delay                 : std_logic      ;
signal fd_main_tm_sech_lw_read_in_progress      : std_logic      ;
signal fd_main_tm_sech_lw_s0                    : std_logic      ;
signal fd_main_tm_sech_lw_s1                    : std_logic      ;
signal fd_main_tm_sech_lw_s2                    : std_logic      ;
signal fd_main_tm_sech_rwsel                    : std_logic      ;
signal fd_main_tm_secl_int_read                 : std_logic_vector(31 downto 0);
signal fd_main_tm_secl_int_write                : std_logic_vector(31 downto 0);
signal fd_main_tm_secl_lw                       : std_logic      ;
signal fd_main_tm_secl_lw_delay                 : std_logic      ;
signal fd_main_tm_secl_lw_read_in_progress      : std_logic      ;
signal fd_main_tm_secl_lw_s0                    : std_logic      ;
signal fd_main_tm_secl_lw_s1                    : std_logic      ;
signal fd_main_tm_secl_lw_s2                    : std_logic      ;
signal fd_main_tm_secl_rwsel                    : std_logic      ;
signal fd_main_tm_cycles_int_read               : std_logic_vector(27 downto 0);
signal fd_main_tm_cycles_int_write              : std_logic_vector(27 downto 0);
signal fd_main_tm_cycles_lw                     : std_logic      ;
signal fd_main_tm_cycles_lw_delay               : std_logic      ;
signal fd_main_tm_cycles_lw_read_in_progress    : std_logic      ;
signal fd_main_tm_cycles_lw_s0                  : std_logic      ;
signal fd_main_tm_cycles_lw_s1                  : std_logic      ;
signal fd_main_tm_cycles_lw_s2                  : std_logic      ;
signal fd_main_tm_cycles_rwsel                  : std_logic      ;
signal fd_main_tdr_int_read                     : std_logic_vector(27 downto 0);
signal fd_main_tdr_int_write                    : std_logic_vector(27 downto 0);
signal fd_main_tdr_lw                           : std_logic      ;
signal fd_main_tdr_lw_delay                     : std_logic      ;
signal fd_main_tdr_lw_read_in_progress          : std_logic      ;
signal fd_main_tdr_lw_s0                        : std_logic      ;
signal fd_main_tdr_lw_s1                        : std_logic      ;
signal fd_main_tdr_lw_s2                        : std_logic      ;
signal fd_main_tdr_rwsel                        : std_logic      ;
signal fd_main_tdcsr_write_int                  : std_logic      ;
signal fd_main_tdcsr_write_int_delay            : std_logic      ;
signal fd_main_tdcsr_write_sync0                : std_logic      ;
signal fd_main_tdcsr_write_sync1                : std_logic      ;
signal fd_main_tdcsr_write_sync2                : std_logic      ;
signal fd_main_tdcsr_read_int                   : std_logic      ;
signal fd_main_tdcsr_read_int_delay             : std_logic      ;
signal fd_main_tdcsr_read_sync0                 : std_logic      ;
signal fd_main_tdcsr_read_sync1                 : std_logic      ;
signal fd_main_tdcsr_read_sync2                 : std_logic      ;
signal fd_main_tdcsr_empty_sync0                : std_logic      ;
signal fd_main_tdcsr_empty_sync1                : std_logic      ;
signal fd_main_tdcsr_stop_en_int                : std_logic      ;
signal fd_main_tdcsr_stop_en_int_delay          : std_logic      ;
signal fd_main_tdcsr_stop_en_sync0              : std_logic      ;
signal fd_main_tdcsr_stop_en_sync1              : std_logic      ;
signal fd_main_tdcsr_stop_en_sync2              : std_logic      ;
signal fd_main_tdcsr_start_dis_int              : std_logic      ;
signal fd_main_tdcsr_start_dis_int_delay        : std_logic      ;
signal fd_main_tdcsr_start_dis_sync0            : std_logic      ;
signal fd_main_tdcsr_start_dis_sync1            : std_logic      ;
signal fd_main_tdcsr_start_dis_sync2            : std_logic      ;
signal fd_main_tdcsr_start_en_int               : std_logic      ;
signal fd_main_tdcsr_start_en_int_delay         : std_logic      ;
signal fd_main_tdcsr_start_en_sync0             : std_logic      ;
signal fd_main_tdcsr_start_en_sync1             : std_logic      ;
signal fd_main_tdcsr_start_en_sync2             : std_logic      ;
signal fd_main_tdcsr_stop_dis_int               : std_logic      ;
signal fd_main_tdcsr_stop_dis_int_delay         : std_logic      ;
signal fd_main_tdcsr_stop_dis_sync0             : std_logic      ;
signal fd_main_tdcsr_stop_dis_sync1             : std_logic      ;
signal fd_main_tdcsr_stop_dis_sync2             : std_logic      ;
signal fd_main_tdcsr_alutrig_int                : std_logic      ;
signal fd_main_tdcsr_alutrig_int_delay          : std_logic      ;
signal fd_main_tdcsr_alutrig_sync0              : std_logic      ;
signal fd_main_tdcsr_alutrig_sync1              : std_logic      ;
signal fd_main_tdcsr_alutrig_sync2              : std_logic      ;
signal fd_main_tdcsr_idelay_ce_int              : std_logic      ;
signal fd_main_tdcsr_idelay_ce_int_delay        : std_logic      ;
signal fd_main_tdcsr_idelay_ce_sync0            : std_logic      ;
signal fd_main_tdcsr_idelay_ce_sync1            : std_logic      ;
signal fd_main_tdcsr_idelay_ce_sync2            : std_logic      ;
signal fd_main_calr_cal_pulse_int               : std_logic      ;
signal fd_main_calr_cal_pulse_int_delay         : std_logic      ;
signal fd_main_calr_cal_pulse_sync0             : std_logic      ;
signal fd_main_calr_cal_pulse_sync1             : std_logic      ;
signal fd_main_calr_cal_pulse_sync2             : std_logic      ;
signal fd_main_calr_cal_pps_int                 : std_logic      ;
signal fd_main_calr_cal_pps_sync0               : std_logic      ;
signal fd_main_calr_cal_pps_sync1               : std_logic      ;
signal fd_main_calr_cal_dmtd_int                : std_logic      ;
signal fd_main_calr_psel_int                    : std_logic_vector(3 downto 0);
signal fd_main_calr_psel_swb                    : std_logic      ;
signal fd_main_calr_psel_swb_delay              : std_logic      ;
signal fd_main_calr_psel_swb_s0                 : std_logic      ;
signal fd_main_calr_psel_swb_s1                 : std_logic      ;
signal fd_main_calr_psel_swb_s2                 : std_logic      ;
signal fd_main_adsfr_int                        : std_logic_vector(17 downto 0);
signal fd_main_adsfr_swb                        : std_logic      ;
signal fd_main_adsfr_swb_delay                  : std_logic      ;
signal fd_main_adsfr_swb_s0                     : std_logic      ;
signal fd_main_adsfr_swb_s1                     : std_logic      ;
signal fd_main_adsfr_swb_s2                     : std_logic      ;
signal fd_main_atmcr_c_thr_int                  : std_logic_vector(7 downto 0);
signal fd_main_atmcr_c_thr_swb                  : std_logic      ;
signal fd_main_atmcr_c_thr_swb_delay            : std_logic      ;
signal fd_main_atmcr_c_thr_swb_s0               : std_logic      ;
signal fd_main_atmcr_c_thr_swb_s1               : std_logic      ;
signal fd_main_atmcr_c_thr_swb_s2               : std_logic      ;
signal fd_main_atmcr_f_thr_int                  : std_logic_vector(22 downto 0);
signal fd_main_atmcr_f_thr_swb                  : std_logic      ;
signal fd_main_atmcr_f_thr_swb_delay            : std_logic      ;
signal fd_main_atmcr_f_thr_swb_s0               : std_logic      ;
signal fd_main_atmcr_f_thr_swb_s1               : std_logic      ;
signal fd_main_atmcr_f_thr_swb_s2               : std_logic      ;
signal fd_main_asor_offset_int                  : std_logic_vector(22 downto 0);
signal fd_main_asor_offset_swb                  : std_logic      ;
signal fd_main_asor_offset_swb_delay            : std_logic      ;
signal fd_main_asor_offset_swb_s0               : std_logic      ;
signal fd_main_asor_offset_swb_s1               : std_logic      ;
signal fd_main_asor_offset_swb_s2               : std_logic      ;
signal fd_main_iecraw_int                       : std_logic_vector(31 downto 0);
signal fd_main_iecraw_lwb                       : std_logic      ;
signal fd_main_iecraw_lwb_delay                 : std_logic      ;
signal fd_main_iecraw_lwb_in_progress           : std_logic      ;
signal fd_main_iecraw_lwb_s0                    : std_logic      ;
signal fd_main_iecraw_lwb_s1                    : std_logic      ;
signal fd_main_iecraw_lwb_s2                    : std_logic      ;
signal fd_main_iectag_int                       : std_logic_vector(31 downto 0);
signal fd_main_iectag_lwb                       : std_logic      ;
signal fd_main_iectag_lwb_delay                 : std_logic      ;
signal fd_main_iectag_lwb_in_progress           : std_logic      ;
signal fd_main_iectag_lwb_s0                    : std_logic      ;
signal fd_main_iectag_lwb_s1                    : std_logic      ;
signal fd_main_iectag_lwb_s2                    : std_logic      ;
signal fd_main_iepd_rst_stat_int                : std_logic      ;
signal fd_main_iepd_rst_stat_int_delay          : std_logic      ;
signal fd_main_iepd_rst_stat_sync0              : std_logic      ;
signal fd_main_iepd_rst_stat_sync1              : std_logic      ;
signal fd_main_iepd_rst_stat_sync2              : std_logic      ;
signal fd_main_iepd_pdelay_int                  : std_logic_vector(7 downto 0);
signal fd_main_iepd_pdelay_lwb                  : std_logic      ;
signal fd_main_iepd_pdelay_lwb_delay            : std_logic      ;
signal fd_main_iepd_pdelay_lwb_in_progress      : std_logic      ;
signal fd_main_iepd_pdelay_lwb_s0               : std_logic      ;
signal fd_main_iepd_pdelay_lwb_s1               : std_logic      ;
signal fd_main_iepd_pdelay_lwb_s2               : std_logic      ;
signal fd_main_scr_sel_dac_int                  : std_logic      ;
signal fd_main_scr_sel_pll_int                  : std_logic      ;
signal fd_main_scr_sel_gpio_int                 : std_logic      ;
signal fd_main_scr_cpol_int                     : std_logic      ;
signal fd_main_scr_start_dly0                   : std_logic      ;
signal fd_main_scr_start_int                    : std_logic      ;
signal fd_main_rcrr_int                         : std_logic_vector(31 downto 0);
signal fd_main_rcrr_lwb                         : std_logic      ;
signal fd_main_rcrr_lwb_delay                   : std_logic      ;
signal fd_main_rcrr_lwb_in_progress             : std_logic      ;
signal fd_main_rcrr_lwb_s0                      : std_logic      ;
signal fd_main_rcrr_lwb_s1                      : std_logic      ;
signal fd_main_rcrr_lwb_s2                      : std_logic      ;
signal fd_main_tsbcr_chan_mask_int              : std_logic_vector(4 downto 0);
signal fd_main_tsbcr_chan_mask_swb              : std_logic      ;
signal fd_main_tsbcr_chan_mask_swb_delay        : std_logic      ;
signal fd_main_tsbcr_chan_mask_swb_s0           : std_logic      ;
signal fd_main_tsbcr_chan_mask_swb_s1           : std_logic      ;
signal fd_main_tsbcr_chan_mask_swb_s2           : std_logic      ;
signal fd_main_tsbcr_enable_int                 : std_logic      ;
signal fd_main_tsbcr_purge_dly0                 : std_logic      ;
signal fd_main_tsbcr_purge_int                  : std_logic      ;
signal fd_main_tsbcr_rst_seq_int                : std_logic      ;
signal fd_main_tsbcr_rst_seq_int_delay          : std_logic      ;
signal fd_main_tsbcr_rst_seq_sync0              : std_logic      ;
signal fd_main_tsbcr_rst_seq_sync1              : std_logic      ;
signal fd_main_tsbcr_rst_seq_sync2              : std_logic      ;
signal fd_main_tsbcr_raw_int                    : std_logic      ;
signal fd_main_tsbir_timeout_int                : std_logic_vector(9 downto 0);
signal fd_main_tsbir_threshold_int              : std_logic_vector(11 downto 0);
signal fd_main_i2cr_scl_out_int                 : std_logic      ;
signal fd_main_i2cr_sda_out_int                 : std_logic      ;
signal fd_main_tder2_pelt_drive_int             : std_logic_vector(31 downto 0);
signal fd_main_tsbr_advance_adv_dly0            : std_logic      ;
signal fd_main_tsbr_advance_adv_int             : std_logic      ;
signal eic_idr_int                              : std_logic_vector(2 downto 0);
signal eic_idr_write_int                        : std_logic      ;
signal eic_ier_int                              : std_logic_vector(2 downto 0);
signal eic_ier_write_int                        : std_logic      ;
signal eic_imr_int                              : std_logic_vector(2 downto 0);
signal eic_isr_clear_int                        : std_logic_vector(2 downto 0);
signal eic_isr_status_int                       : std_logic_vector(2 downto 0);
signal eic_irq_ack_int                          : std_logic_vector(2 downto 0);
signal eic_isr_write_int                        : std_logic      ;
signal irq_inputs_vector_int                    : std_logic_vector(2 downto 0);
signal ack_sreg                                 : std_logic_vector(9 downto 0);
signal rddata_reg                               : std_logic_vector(31 downto 0);
signal wrdata_reg                               : std_logic_vector(31 downto 0);
signal bwsel_reg                                : std_logic_vector(3 downto 0);
signal rwaddr_reg                               : std_logic_vector(5 downto 0);
signal ack_in_progress                          : std_logic      ;
signal wr_int                                   : std_logic      ;
signal rd_int                                   : std_logic      ;
signal allones                                  : std_logic_vector(31 downto 0);
signal allzeros                                 : std_logic_vector(31 downto 0);

begin
-- Some internal signals assignments
wrdata_reg <= wb_dat_i;
-- 
-- Main register bank access process.
process (clk_sys_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    ack_sreg <= "0000000000";
    ack_in_progress <= '0';
    rddata_reg <= "00000000000000000000000000000000";
    regs_o.rstr_rst_fmc_wr_o <= '0';
    regs_o.rstr_rst_core_wr_o <= '0';
    regs_o.rstr_lock_wr_o <= '0';
    fd_main_gcr_bypass_int <= '0';
    fd_main_gcr_input_en_int <= '0';
    tcr_rd_ack_o <= '0';
    fd_main_tcr_wr_enable_int <= '0';
    fd_main_tcr_cap_time_int <= '0';
    fd_main_tcr_cap_time_int_delay <= '0';
    fd_main_tcr_set_time_int <= '0';
    fd_main_tcr_set_time_int_delay <= '0';
    fd_main_tm_sech_lw <= '0';
    fd_main_tm_sech_lw_delay <= '0';
    fd_main_tm_sech_lw_read_in_progress <= '0';
    fd_main_tm_sech_rwsel <= '0';
    fd_main_tm_sech_int_write <= "00000000";
    fd_main_tm_secl_lw <= '0';
    fd_main_tm_secl_lw_delay <= '0';
    fd_main_tm_secl_lw_read_in_progress <= '0';
    fd_main_tm_secl_rwsel <= '0';
    fd_main_tm_secl_int_write <= "00000000000000000000000000000000";
    fd_main_tm_cycles_lw <= '0';
    fd_main_tm_cycles_lw_delay <= '0';
    fd_main_tm_cycles_lw_read_in_progress <= '0';
    fd_main_tm_cycles_rwsel <= '0';
    fd_main_tm_cycles_int_write <= "0000000000000000000000000000";
    fd_main_tdr_lw <= '0';
    fd_main_tdr_lw_delay <= '0';
    fd_main_tdr_lw_read_in_progress <= '0';
    fd_main_tdr_rwsel <= '0';
    fd_main_tdr_int_write <= "0000000000000000000000000000";
    fd_main_tdcsr_write_int <= '0';
    fd_main_tdcsr_write_int_delay <= '0';
    fd_main_tdcsr_read_int <= '0';
    fd_main_tdcsr_read_int_delay <= '0';
    fd_main_tdcsr_stop_en_int <= '0';
    fd_main_tdcsr_stop_en_int_delay <= '0';
    fd_main_tdcsr_start_dis_int <= '0';
    fd_main_tdcsr_start_dis_int_delay <= '0';
    fd_main_tdcsr_start_en_int <= '0';
    fd_main_tdcsr_start_en_int_delay <= '0';
    fd_main_tdcsr_stop_dis_int <= '0';
    fd_main_tdcsr_stop_dis_int_delay <= '0';
    fd_main_tdcsr_alutrig_int <= '0';
    fd_main_tdcsr_alutrig_int_delay <= '0';
    fd_main_tdcsr_idelay_ce_int <= '0';
    fd_main_tdcsr_idelay_ce_int_delay <= '0';
    fd_main_calr_cal_pulse_int <= '0';
    fd_main_calr_cal_pulse_int_delay <= '0';
    fd_main_calr_cal_pps_int <= '0';
    fd_main_calr_cal_dmtd_int <= '0';
    fd_main_calr_psel_int <= "0000";
    fd_main_calr_psel_swb <= '0';
    fd_main_calr_psel_swb_delay <= '0';
    dmtr_in_rd_ack_o <= '0';
    dmtr_out_rd_ack_o <= '0';
    fd_main_adsfr_int <= "000000000000000000";
    fd_main_adsfr_swb <= '0';
    fd_main_adsfr_swb_delay <= '0';
    fd_main_atmcr_c_thr_int <= "00000000";
    fd_main_atmcr_c_thr_swb <= '0';
    fd_main_atmcr_c_thr_swb_delay <= '0';
    fd_main_atmcr_f_thr_int <= "00000000000000000000000";
    fd_main_atmcr_f_thr_swb <= '0';
    fd_main_atmcr_f_thr_swb_delay <= '0';
    fd_main_asor_offset_int <= "00000000000000000000000";
    fd_main_asor_offset_swb <= '0';
    fd_main_asor_offset_swb_delay <= '0';
    fd_main_iecraw_lwb <= '0';
    fd_main_iecraw_lwb_delay <= '0';
    fd_main_iecraw_lwb_in_progress <= '0';
    fd_main_iectag_lwb <= '0';
    fd_main_iectag_lwb_delay <= '0';
    fd_main_iectag_lwb_in_progress <= '0';
    fd_main_iepd_rst_stat_int <= '0';
    fd_main_iepd_rst_stat_int_delay <= '0';
    fd_main_iepd_pdelay_lwb <= '0';
    fd_main_iepd_pdelay_lwb_delay <= '0';
    fd_main_iepd_pdelay_lwb_in_progress <= '0';
    regs_o.scr_data_load_o <= '0';
    fd_main_scr_sel_dac_int <= '0';
    fd_main_scr_sel_pll_int <= '0';
    fd_main_scr_sel_gpio_int <= '0';
    fd_main_scr_cpol_int <= '0';
    fd_main_scr_start_int <= '0';
    fd_main_rcrr_lwb <= '0';
    fd_main_rcrr_lwb_delay <= '0';
    fd_main_rcrr_lwb_in_progress <= '0';
    fd_main_tsbcr_chan_mask_int <= "00000";
    fd_main_tsbcr_chan_mask_swb <= '0';
    fd_main_tsbcr_chan_mask_swb_delay <= '0';
    fd_main_tsbcr_enable_int <= '0';
    fd_main_tsbcr_purge_int <= '0';
    fd_main_tsbcr_rst_seq_int <= '0';
    fd_main_tsbcr_rst_seq_int_delay <= '0';
    tsbcr_read_ack_o <= '0';
    fd_main_tsbcr_raw_int <= '0';
    fd_main_tsbir_timeout_int <= "0000000000";
    fd_main_tsbir_threshold_int <= "000000000000";
    fid_read_ack_o <= '0';
    fd_main_i2cr_scl_out_int <= '1';
    fd_main_i2cr_sda_out_int <= '1';
    fd_main_tder2_pelt_drive_int <= "00000000000000000000000000000000";
    fd_main_tsbr_advance_adv_int <= '0';
    regs_o.iodelay_adj_n_taps_load_o <= '0';
    eic_idr_write_int <= '0';
    eic_ier_write_int <= '0';
    eic_isr_write_int <= '0';
  elsif rising_edge(clk_sys_i) then
-- advance the ACK generator shift register
    ack_sreg(8 downto 0) <= ack_sreg(9 downto 1);
    ack_sreg(9) <= '0';
    if (ack_in_progress = '1') then
      if (ack_sreg(0) = '1') then
        regs_o.rstr_rst_fmc_wr_o <= '0';
        regs_o.rstr_rst_core_wr_o <= '0';
        regs_o.rstr_lock_wr_o <= '0';
        tcr_rd_ack_o <= '0';
        dmtr_in_rd_ack_o <= '0';
        dmtr_out_rd_ack_o <= '0';
        regs_o.scr_data_load_o <= '0';
        fd_main_scr_start_int <= '0';
        fd_main_tsbcr_purge_int <= '0';
        tsbcr_read_ack_o <= '0';
        fid_read_ack_o <= '0';
        fd_main_tsbr_advance_adv_int <= '0';
        regs_o.iodelay_adj_n_taps_load_o <= '0';
        eic_idr_write_int <= '0';
        eic_ier_write_int <= '0';
        eic_isr_write_int <= '0';
        ack_in_progress <= '0';
      else
        regs_o.rstr_rst_fmc_wr_o <= '0';
        regs_o.rstr_rst_core_wr_o <= '0';
        regs_o.rstr_lock_wr_o <= '0';
        fd_main_tcr_cap_time_int <= fd_main_tcr_cap_time_int_delay;
        fd_main_tcr_cap_time_int_delay <= '0';
        fd_main_tcr_set_time_int <= fd_main_tcr_set_time_int_delay;
        fd_main_tcr_set_time_int_delay <= '0';
        fd_main_tm_sech_lw <= fd_main_tm_sech_lw_delay;
        fd_main_tm_sech_lw_delay <= '0';
        if ((ack_sreg(1) = '1') and (fd_main_tm_sech_lw_read_in_progress = '1')) then
          rddata_reg(7 downto 0) <= fd_main_tm_sech_int_read;
          fd_main_tm_sech_lw_read_in_progress <= '0';
        end if;
        fd_main_tm_secl_lw <= fd_main_tm_secl_lw_delay;
        fd_main_tm_secl_lw_delay <= '0';
        if ((ack_sreg(1) = '1') and (fd_main_tm_secl_lw_read_in_progress = '1')) then
          rddata_reg(31 downto 0) <= fd_main_tm_secl_int_read;
          fd_main_tm_secl_lw_read_in_progress <= '0';
        end if;
        fd_main_tm_cycles_lw <= fd_main_tm_cycles_lw_delay;
        fd_main_tm_cycles_lw_delay <= '0';
        if ((ack_sreg(1) = '1') and (fd_main_tm_cycles_lw_read_in_progress = '1')) then
          rddata_reg(27 downto 0) <= fd_main_tm_cycles_int_read;
          fd_main_tm_cycles_lw_read_in_progress <= '0';
        end if;
        fd_main_tdr_lw <= fd_main_tdr_lw_delay;
        fd_main_tdr_lw_delay <= '0';
        if ((ack_sreg(1) = '1') and (fd_main_tdr_lw_read_in_progress = '1')) then
          rddata_reg(27 downto 0) <= fd_main_tdr_int_read;
          fd_main_tdr_lw_read_in_progress <= '0';
        end if;
        fd_main_tdcsr_write_int <= fd_main_tdcsr_write_int_delay;
        fd_main_tdcsr_write_int_delay <= '0';
        fd_main_tdcsr_read_int <= fd_main_tdcsr_read_int_delay;
        fd_main_tdcsr_read_int_delay <= '0';
        fd_main_tdcsr_stop_en_int <= fd_main_tdcsr_stop_en_int_delay;
        fd_main_tdcsr_stop_en_int_delay <= '0';
        fd_main_tdcsr_start_dis_int <= fd_main_tdcsr_start_dis_int_delay;
        fd_main_tdcsr_start_dis_int_delay <= '0';
        fd_main_tdcsr_start_en_int <= fd_main_tdcsr_start_en_int_delay;
        fd_main_tdcsr_start_en_int_delay <= '0';
        fd_main_tdcsr_stop_dis_int <= fd_main_tdcsr_stop_dis_int_delay;
        fd_main_tdcsr_stop_dis_int_delay <= '0';
        fd_main_tdcsr_alutrig_int <= fd_main_tdcsr_alutrig_int_delay;
        fd_main_tdcsr_alutrig_int_delay <= '0';
        fd_main_tdcsr_idelay_ce_int <= fd_main_tdcsr_idelay_ce_int_delay;
        fd_main_tdcsr_idelay_ce_int_delay <= '0';
        fd_main_calr_cal_pulse_int <= fd_main_calr_cal_pulse_int_delay;
        fd_main_calr_cal_pulse_int_delay <= '0';
        fd_main_calr_psel_swb <= fd_main_calr_psel_swb_delay;
        fd_main_calr_psel_swb_delay <= '0';
        fd_main_adsfr_swb <= fd_main_adsfr_swb_delay;
        fd_main_adsfr_swb_delay <= '0';
        fd_main_atmcr_c_thr_swb <= fd_main_atmcr_c_thr_swb_delay;
        fd_main_atmcr_c_thr_swb_delay <= '0';
        fd_main_atmcr_f_thr_swb <= fd_main_atmcr_f_thr_swb_delay;
        fd_main_atmcr_f_thr_swb_delay <= '0';
        fd_main_asor_offset_swb <= fd_main_asor_offset_swb_delay;
        fd_main_asor_offset_swb_delay <= '0';
        fd_main_iecraw_lwb <= fd_main_iecraw_lwb_delay;
        fd_main_iecraw_lwb_delay <= '0';
        if ((ack_sreg(1) = '1') and (fd_main_iecraw_lwb_in_progress = '1')) then
          rddata_reg(31 downto 0) <= fd_main_iecraw_int;
          fd_main_iecraw_lwb_in_progress <= '0';
        end if;
        fd_main_iectag_lwb <= fd_main_iectag_lwb_delay;
        fd_main_iectag_lwb_delay <= '0';
        if ((ack_sreg(1) = '1') and (fd_main_iectag_lwb_in_progress = '1')) then
          rddata_reg(31 downto 0) <= fd_main_iectag_int;
          fd_main_iectag_lwb_in_progress <= '0';
        end if;
        fd_main_iepd_rst_stat_int <= fd_main_iepd_rst_stat_int_delay;
        fd_main_iepd_rst_stat_int_delay <= '0';
        fd_main_iepd_pdelay_lwb <= fd_main_iepd_pdelay_lwb_delay;
        fd_main_iepd_pdelay_lwb_delay <= '0';
        if ((ack_sreg(1) = '1') and (fd_main_iepd_pdelay_lwb_in_progress = '1')) then
          rddata_reg(8 downto 1) <= fd_main_iepd_pdelay_int;
          fd_main_iepd_pdelay_lwb_in_progress <= '0';
        end if;
        regs_o.scr_data_load_o <= '0';
        fd_main_rcrr_lwb <= fd_main_rcrr_lwb_delay;
        fd_main_rcrr_lwb_delay <= '0';
        if ((ack_sreg(1) = '1') and (fd_main_rcrr_lwb_in_progress = '1')) then
          rddata_reg(31 downto 0) <= fd_main_rcrr_int;
          fd_main_rcrr_lwb_in_progress <= '0';
        end if;
        fd_main_tsbcr_chan_mask_swb <= fd_main_tsbcr_chan_mask_swb_delay;
        fd_main_tsbcr_chan_mask_swb_delay <= '0';
        fd_main_tsbcr_rst_seq_int <= fd_main_tsbcr_rst_seq_int_delay;
        fd_main_tsbcr_rst_seq_int_delay <= '0';
        regs_o.iodelay_adj_n_taps_load_o <= '0';
      end if;
    else
      if ((wb_cyc_i = '1') and (wb_stb_i = '1')) then
        case rwaddr_reg(5 downto 0) is
        when "000000" => 
          if (wb_we_i = '1') then
            regs_o.rstr_rst_fmc_wr_o <= '1';
            regs_o.rstr_rst_core_wr_o <= '1';
            regs_o.rstr_lock_wr_o <= '1';
          end if;
          rddata_reg(0) <= 'X';
          rddata_reg(1) <= 'X';
          rddata_reg(2) <= 'X';
          rddata_reg(3) <= 'X';
          rddata_reg(4) <= 'X';
          rddata_reg(5) <= 'X';
          rddata_reg(6) <= 'X';
          rddata_reg(7) <= 'X';
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "000001" => 
          if (wb_we_i = '1') then
          end if;
          rddata_reg(31 downto 0) <= "11110001100111101101111000011010";
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "000010" => 
          if (wb_we_i = '1') then
            fd_main_gcr_bypass_int <= wrdata_reg(0);
            fd_main_gcr_input_en_int <= wrdata_reg(1);
          end if;
          rddata_reg(0) <= fd_main_gcr_bypass_int;
          rddata_reg(1) <= fd_main_gcr_input_en_int;
          rddata_reg(2) <= regs_i.gcr_ddr_locked_i;
          rddata_reg(3) <= regs_i.gcr_fmc_present_i;
          rddata_reg(4) <= 'X';
          rddata_reg(5) <= 'X';
          rddata_reg(6) <= 'X';
          rddata_reg(7) <= 'X';
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(3) <= '1';
          ack_in_progress <= '1';
        when "000011" => 
          if (wb_we_i = '1') then
            fd_main_tcr_wr_enable_int <= wrdata_reg(1);
            fd_main_tcr_cap_time_int <= wrdata_reg(6);
            fd_main_tcr_cap_time_int_delay <= wrdata_reg(6);
            fd_main_tcr_set_time_int <= wrdata_reg(7);
            fd_main_tcr_set_time_int_delay <= wrdata_reg(7);
          end if;
          rddata_reg(0) <= regs_i.tcr_dmtd_stat_i;
          tcr_rd_ack_o <= '1';
          rddata_reg(1) <= fd_main_tcr_wr_enable_int;
          rddata_reg(2) <= regs_i.tcr_wr_locked_i;
          rddata_reg(3) <= regs_i.tcr_wr_present_i;
          rddata_reg(4) <= regs_i.tcr_wr_ready_i;
          rddata_reg(5) <= regs_i.tcr_wr_link_i;
          rddata_reg(6) <= '0';
          rddata_reg(7) <= '0';
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(4) <= '1';
          ack_in_progress <= '1';
        when "000100" => 
          if (wb_we_i = '1') then
            fd_main_tm_sech_int_write <= wrdata_reg(7 downto 0);
            fd_main_tm_sech_lw <= '1';
            fd_main_tm_sech_lw_delay <= '1';
            fd_main_tm_sech_lw_read_in_progress <= '0';
            fd_main_tm_sech_rwsel <= '1';
          end if;
          if (wb_we_i = '0') then
            fd_main_tm_sech_lw <= '1';
            fd_main_tm_sech_lw_delay <= '1';
            fd_main_tm_sech_lw_read_in_progress <= '1';
            fd_main_tm_sech_rwsel <= '0';
          end if;
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(5) <= '1';
          ack_in_progress <= '1';
        when "000101" => 
          if (wb_we_i = '1') then
            fd_main_tm_secl_int_write <= wrdata_reg(31 downto 0);
            fd_main_tm_secl_lw <= '1';
            fd_main_tm_secl_lw_delay <= '1';
            fd_main_tm_secl_lw_read_in_progress <= '0';
            fd_main_tm_secl_rwsel <= '1';
          end if;
          if (wb_we_i = '0') then
            fd_main_tm_secl_lw <= '1';
            fd_main_tm_secl_lw_delay <= '1';
            fd_main_tm_secl_lw_read_in_progress <= '1';
            fd_main_tm_secl_rwsel <= '0';
          end if;
          ack_sreg(5) <= '1';
          ack_in_progress <= '1';
        when "000110" => 
          if (wb_we_i = '1') then
            fd_main_tm_cycles_int_write <= wrdata_reg(27 downto 0);
            fd_main_tm_cycles_lw <= '1';
            fd_main_tm_cycles_lw_delay <= '1';
            fd_main_tm_cycles_lw_read_in_progress <= '0';
            fd_main_tm_cycles_rwsel <= '1';
          end if;
          if (wb_we_i = '0') then
            fd_main_tm_cycles_lw <= '1';
            fd_main_tm_cycles_lw_delay <= '1';
            fd_main_tm_cycles_lw_read_in_progress <= '1';
            fd_main_tm_cycles_rwsel <= '0';
          end if;
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(5) <= '1';
          ack_in_progress <= '1';
        when "000111" => 
          if (wb_we_i = '1') then
            fd_main_tdr_int_write <= wrdata_reg(27 downto 0);
            fd_main_tdr_lw <= '1';
            fd_main_tdr_lw_delay <= '1';
            fd_main_tdr_lw_read_in_progress <= '0';
            fd_main_tdr_rwsel <= '1';
          end if;
          if (wb_we_i = '0') then
            fd_main_tdr_lw <= '1';
            fd_main_tdr_lw_delay <= '1';
            fd_main_tdr_lw_read_in_progress <= '1';
            fd_main_tdr_rwsel <= '0';
          end if;
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(5) <= '1';
          ack_in_progress <= '1';
        when "001000" => 
          if (wb_we_i = '1') then
            fd_main_tdcsr_write_int <= wrdata_reg(0);
            fd_main_tdcsr_write_int_delay <= wrdata_reg(0);
            fd_main_tdcsr_read_int <= wrdata_reg(1);
            fd_main_tdcsr_read_int_delay <= wrdata_reg(1);
            fd_main_tdcsr_stop_en_int <= wrdata_reg(3);
            fd_main_tdcsr_stop_en_int_delay <= wrdata_reg(3);
            fd_main_tdcsr_start_dis_int <= wrdata_reg(4);
            fd_main_tdcsr_start_dis_int_delay <= wrdata_reg(4);
            fd_main_tdcsr_start_en_int <= wrdata_reg(5);
            fd_main_tdcsr_start_en_int_delay <= wrdata_reg(5);
            fd_main_tdcsr_stop_dis_int <= wrdata_reg(6);
            fd_main_tdcsr_stop_dis_int_delay <= wrdata_reg(6);
            fd_main_tdcsr_alutrig_int <= wrdata_reg(7);
            fd_main_tdcsr_alutrig_int_delay <= wrdata_reg(7);
            fd_main_tdcsr_idelay_ce_int <= wrdata_reg(8);
            fd_main_tdcsr_idelay_ce_int_delay <= wrdata_reg(8);
          end if;
          rddata_reg(0) <= '0';
          rddata_reg(1) <= '0';
          rddata_reg(2) <= fd_main_tdcsr_empty_sync1;
          rddata_reg(3) <= '0';
          rddata_reg(4) <= '0';
          rddata_reg(5) <= '0';
          rddata_reg(6) <= '0';
          rddata_reg(7) <= '0';
          rddata_reg(8) <= '0';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(4) <= '1';
          ack_in_progress <= '1';
        when "001001" => 
          if (wb_we_i = '1') then
            fd_main_calr_cal_pulse_int <= wrdata_reg(0);
            fd_main_calr_cal_pulse_int_delay <= wrdata_reg(0);
            fd_main_calr_cal_pps_int <= wrdata_reg(1);
            fd_main_calr_cal_dmtd_int <= wrdata_reg(2);
            fd_main_calr_psel_int <= wrdata_reg(6 downto 3);
            fd_main_calr_psel_swb <= '1';
            fd_main_calr_psel_swb_delay <= '1';
          end if;
          rddata_reg(0) <= '0';
          rddata_reg(1) <= fd_main_calr_cal_pps_int;
          rddata_reg(2) <= fd_main_calr_cal_dmtd_int;
          rddata_reg(6 downto 3) <= fd_main_calr_psel_int;
          rddata_reg(7) <= 'X';
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(4) <= '1';
          ack_in_progress <= '1';
        when "001010" => 
          if (wb_we_i = '1') then
          end if;
          rddata_reg(30 downto 0) <= regs_i.dmtr_in_tag_i;
          dmtr_in_rd_ack_o <= '1';
          rddata_reg(31) <= regs_i.dmtr_in_rdy_i;
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "001011" => 
          if (wb_we_i = '1') then
          end if;
          rddata_reg(30 downto 0) <= regs_i.dmtr_out_tag_i;
          dmtr_out_rd_ack_o <= '1';
          rddata_reg(31) <= regs_i.dmtr_out_rdy_i;
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "001100" => 
          if (wb_we_i = '1') then
            fd_main_adsfr_int <= wrdata_reg(17 downto 0);
            fd_main_adsfr_swb <= '1';
            fd_main_adsfr_swb_delay <= '1';
          end if;
          rddata_reg(17 downto 0) <= fd_main_adsfr_int;
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(3) <= '1';
          ack_in_progress <= '1';
        when "001101" => 
          if (wb_we_i = '1') then
            fd_main_atmcr_c_thr_int <= wrdata_reg(7 downto 0);
            fd_main_atmcr_c_thr_swb <= '1';
            fd_main_atmcr_c_thr_swb_delay <= '1';
            fd_main_atmcr_f_thr_int <= wrdata_reg(30 downto 8);
            fd_main_atmcr_f_thr_swb <= '1';
            fd_main_atmcr_f_thr_swb_delay <= '1';
          end if;
          rddata_reg(7 downto 0) <= fd_main_atmcr_c_thr_int;
          rddata_reg(30 downto 8) <= fd_main_atmcr_f_thr_int;
          rddata_reg(31) <= 'X';
          ack_sreg(3) <= '1';
          ack_in_progress <= '1';
        when "001110" => 
          if (wb_we_i = '1') then
            fd_main_asor_offset_int <= wrdata_reg(22 downto 0);
            fd_main_asor_offset_swb <= '1';
            fd_main_asor_offset_swb_delay <= '1';
          end if;
          rddata_reg(22 downto 0) <= fd_main_asor_offset_int;
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(3) <= '1';
          ack_in_progress <= '1';
        when "001111" => 
          if (wb_we_i = '1') then
          end if;
          if (wb_we_i = '0') then
            fd_main_iecraw_lwb <= '1';
            fd_main_iecraw_lwb_delay <= '1';
            fd_main_iecraw_lwb_in_progress <= '1';
          end if;
          ack_sreg(5) <= '1';
          ack_in_progress <= '1';
        when "010000" => 
          if (wb_we_i = '1') then
          end if;
          if (wb_we_i = '0') then
            fd_main_iectag_lwb <= '1';
            fd_main_iectag_lwb_delay <= '1';
            fd_main_iectag_lwb_in_progress <= '1';
          end if;
          ack_sreg(5) <= '1';
          ack_in_progress <= '1';
        when "010001" => 
          if (wb_we_i = '1') then
            fd_main_iepd_rst_stat_int <= wrdata_reg(0);
            fd_main_iepd_rst_stat_int_delay <= wrdata_reg(0);
          end if;
          rddata_reg(0) <= '0';
          if (wb_we_i = '0') then
            fd_main_iepd_pdelay_lwb <= '1';
            fd_main_iepd_pdelay_lwb_delay <= '1';
            fd_main_iepd_pdelay_lwb_in_progress <= '1';
          end if;
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(5) <= '1';
          ack_in_progress <= '1';
        when "010010" => 
          if (wb_we_i = '1') then
            regs_o.scr_data_load_o <= '1';
            fd_main_scr_sel_dac_int <= wrdata_reg(24);
            fd_main_scr_sel_pll_int <= wrdata_reg(25);
            fd_main_scr_sel_gpio_int <= wrdata_reg(26);
            fd_main_scr_cpol_int <= wrdata_reg(28);
            fd_main_scr_start_int <= wrdata_reg(29);
          end if;
          rddata_reg(23 downto 0) <= regs_i.scr_data_i;
          rddata_reg(24) <= fd_main_scr_sel_dac_int;
          rddata_reg(25) <= fd_main_scr_sel_pll_int;
          rddata_reg(26) <= fd_main_scr_sel_gpio_int;
          rddata_reg(27) <= regs_i.scr_ready_i;
          rddata_reg(28) <= fd_main_scr_cpol_int;
          rddata_reg(29) <= '0';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(2) <= '1';
          ack_in_progress <= '1';
        when "010011" => 
          if (wb_we_i = '1') then
          end if;
          if (wb_we_i = '0') then
            fd_main_rcrr_lwb <= '1';
            fd_main_rcrr_lwb_delay <= '1';
            fd_main_rcrr_lwb_in_progress <= '1';
          end if;
          ack_sreg(5) <= '1';
          ack_in_progress <= '1';
        when "010100" => 
          if (wb_we_i = '1') then
            fd_main_tsbcr_chan_mask_int <= wrdata_reg(4 downto 0);
            fd_main_tsbcr_chan_mask_swb <= '1';
            fd_main_tsbcr_chan_mask_swb_delay <= '1';
            fd_main_tsbcr_enable_int <= wrdata_reg(5);
            fd_main_tsbcr_purge_int <= wrdata_reg(6);
            fd_main_tsbcr_rst_seq_int <= wrdata_reg(7);
            fd_main_tsbcr_rst_seq_int_delay <= wrdata_reg(7);
            fd_main_tsbcr_raw_int <= wrdata_reg(22);
          end if;
          rddata_reg(4 downto 0) <= fd_main_tsbcr_chan_mask_int;
          rddata_reg(5) <= fd_main_tsbcr_enable_int;
          rddata_reg(6) <= '0';
          rddata_reg(7) <= '0';
          rddata_reg(8) <= regs_i.tsbcr_full_i;
          rddata_reg(9) <= regs_i.tsbcr_empty_i;
          tsbcr_read_ack_o <= '1';
          rddata_reg(21 downto 10) <= regs_i.tsbcr_count_i;
          rddata_reg(22) <= fd_main_tsbcr_raw_int;
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(4) <= '1';
          ack_in_progress <= '1';
        when "010101" => 
          if (wb_we_i = '1') then
            fd_main_tsbir_timeout_int <= wrdata_reg(9 downto 0);
            fd_main_tsbir_threshold_int <= wrdata_reg(21 downto 10);
          end if;
          rddata_reg(9 downto 0) <= fd_main_tsbir_timeout_int;
          rddata_reg(21 downto 10) <= fd_main_tsbir_threshold_int;
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "010110" => 
          if (wb_we_i = '1') then
          end if;
          rddata_reg(7 downto 0) <= regs_i.tsbr_sech_i;
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "010111" => 
          if (wb_we_i = '1') then
          end if;
          rddata_reg(31 downto 0) <= regs_i.tsbr_secl_i;
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "011000" => 
          if (wb_we_i = '1') then
          end if;
          rddata_reg(27 downto 0) <= regs_i.tsbr_cycles_i;
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "011001" => 
          if (wb_we_i = '1') then
          end if;
          rddata_reg(3 downto 0) <= regs_i.tsbr_fid_channel_i;
          rddata_reg(15 downto 4) <= regs_i.tsbr_fid_fine_i;
          rddata_reg(31 downto 16) <= regs_i.tsbr_fid_seqid_i;
          fid_read_ack_o <= '1';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "011010" => 
          if (wb_we_i = '1') then
            fd_main_i2cr_scl_out_int <= wrdata_reg(0);
            fd_main_i2cr_sda_out_int <= wrdata_reg(1);
          end if;
          rddata_reg(0) <= fd_main_i2cr_scl_out_int;
          rddata_reg(1) <= fd_main_i2cr_sda_out_int;
          rddata_reg(2) <= regs_i.i2cr_scl_in_i;
          rddata_reg(3) <= regs_i.i2cr_sda_in_i;
          rddata_reg(4) <= 'X';
          rddata_reg(5) <= 'X';
          rddata_reg(6) <= 'X';
          rddata_reg(7) <= 'X';
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "011011" => 
          if (wb_we_i = '1') then
          end if;
          rddata_reg(31 downto 0) <= regs_i.tder1_vcxo_freq_i;
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "011100" => 
          if (wb_we_i = '1') then
            fd_main_tder2_pelt_drive_int <= wrdata_reg(31 downto 0);
          end if;
          rddata_reg(31 downto 0) <= fd_main_tder2_pelt_drive_int;
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "011101" => 
          if (wb_we_i = '1') then
          end if;
          rddata_reg(31 downto 0) <= regs_i.tsbr_debug_i;
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "011110" => 
          if (wb_we_i = '1') then
            fd_main_tsbr_advance_adv_int <= wrdata_reg(0);
          end if;
          rddata_reg(0) <= '0';
          rddata_reg(0) <= 'X';
          rddata_reg(1) <= 'X';
          rddata_reg(2) <= 'X';
          rddata_reg(3) <= 'X';
          rddata_reg(4) <= 'X';
          rddata_reg(5) <= 'X';
          rddata_reg(6) <= 'X';
          rddata_reg(7) <= 'X';
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(2) <= '1';
          ack_in_progress <= '1';
        when "011111" => 
          if (wb_we_i = '1') then
          end if;
          rddata_reg(3 downto 0) <= regs_i.fmc_slot_id_slot_id_i;
          rddata_reg(4) <= 'X';
          rddata_reg(5) <= 'X';
          rddata_reg(6) <= 'X';
          rddata_reg(7) <= 'X';
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "100000" => 
          if (wb_we_i = '1') then
            regs_o.iodelay_adj_n_taps_load_o <= '1';
          end if;
          rddata_reg(7 downto 0) <= regs_i.iodelay_adj_n_taps_i;
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "101000" => 
          if (wb_we_i = '1') then
            eic_idr_write_int <= '1';
          end if;
          rddata_reg(0) <= 'X';
          rddata_reg(1) <= 'X';
          rddata_reg(2) <= 'X';
          rddata_reg(3) <= 'X';
          rddata_reg(4) <= 'X';
          rddata_reg(5) <= 'X';
          rddata_reg(6) <= 'X';
          rddata_reg(7) <= 'X';
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "101001" => 
          if (wb_we_i = '1') then
            eic_ier_write_int <= '1';
          end if;
          rddata_reg(0) <= 'X';
          rddata_reg(1) <= 'X';
          rddata_reg(2) <= 'X';
          rddata_reg(3) <= 'X';
          rddata_reg(4) <= 'X';
          rddata_reg(5) <= 'X';
          rddata_reg(6) <= 'X';
          rddata_reg(7) <= 'X';
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "101010" => 
          if (wb_we_i = '1') then
          end if;
          rddata_reg(2 downto 0) <= eic_imr_int(2 downto 0);
          rddata_reg(3) <= 'X';
          rddata_reg(4) <= 'X';
          rddata_reg(5) <= 'X';
          rddata_reg(6) <= 'X';
          rddata_reg(7) <= 'X';
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "101011" => 
          if (wb_we_i = '1') then
            eic_isr_write_int <= '1';
          end if;
          rddata_reg(2 downto 0) <= eic_isr_status_int(2 downto 0);
          rddata_reg(3) <= 'X';
          rddata_reg(4) <= 'X';
          rddata_reg(5) <= 'X';
          rddata_reg(6) <= 'X';
          rddata_reg(7) <= 'X';
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when others =>
-- prevent the slave from hanging the bus on invalid address
          ack_in_progress <= '1';
          ack_sreg(0) <= '1';
        end case;
      end if;
    end if;
  end if;
end process;


-- Drive the data output bus
wb_dat_o <= rddata_reg;
-- State of the reset Line of the Mezzanine (EXT_RST_N pin)
-- pass-through field: State of the reset Line of the Mezzanine (EXT_RST_N pin) in register: Reset Register
regs_o.rstr_rst_fmc_o <= wrdata_reg(0);
-- State of the reset of the Fine Delay Core
-- pass-through field: State of the reset of the Fine Delay Core in register: Reset Register
regs_o.rstr_rst_core_o <= wrdata_reg(1);
-- Reset magic value
-- pass-through field: Reset magic value in register: Reset Register
regs_o.rstr_lock_o <= wrdata_reg(31 downto 16);
-- Bypass hardware TDC controller
-- synchronizer chain for field : Bypass hardware TDC controller (type RW/RO, clk_sys_i <-> clk_ref_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.gcr_bypass_o <= '0';
    fd_main_gcr_bypass_sync0 <= '0';
    fd_main_gcr_bypass_sync1 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_gcr_bypass_sync0 <= fd_main_gcr_bypass_int;
    fd_main_gcr_bypass_sync1 <= fd_main_gcr_bypass_sync0;
    regs_o.gcr_bypass_o <= fd_main_gcr_bypass_sync1;
  end if;
end process;


-- Enable trigger input
-- synchronizer chain for field : Enable trigger input (type RW/RO, clk_sys_i <-> clk_ref_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.gcr_input_en_o <= '0';
    fd_main_gcr_input_en_sync0 <= '0';
    fd_main_gcr_input_en_sync1 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_gcr_input_en_sync0 <= fd_main_gcr_input_en_int;
    fd_main_gcr_input_en_sync1 <= fd_main_gcr_input_en_sync0;
    regs_o.gcr_input_en_o <= fd_main_gcr_input_en_sync1;
  end if;
end process;


-- PLL lock status
-- Mezzanine present
-- DMTD Clock Status
-- WR Timing Enable
regs_o.tcr_wr_enable_o <= fd_main_tcr_wr_enable_int;
-- WR Timing Locked
-- WR Core Present
-- WR Core Time Ready
-- WR Core Link Up
-- Capture Current Time
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.tcr_cap_time_o <= '0';
    fd_main_tcr_cap_time_sync0 <= '0';
    fd_main_tcr_cap_time_sync1 <= '0';
    fd_main_tcr_cap_time_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_tcr_cap_time_sync0 <= fd_main_tcr_cap_time_int;
    fd_main_tcr_cap_time_sync1 <= fd_main_tcr_cap_time_sync0;
    fd_main_tcr_cap_time_sync2 <= fd_main_tcr_cap_time_sync1;
    regs_o.tcr_cap_time_o <= fd_main_tcr_cap_time_sync2 and (not fd_main_tcr_cap_time_sync1);
  end if;
end process;


-- Set Current Time
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.tcr_set_time_o <= '0';
    fd_main_tcr_set_time_sync0 <= '0';
    fd_main_tcr_set_time_sync1 <= '0';
    fd_main_tcr_set_time_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_tcr_set_time_sync0 <= fd_main_tcr_set_time_int;
    fd_main_tcr_set_time_sync1 <= fd_main_tcr_set_time_sync0;
    fd_main_tcr_set_time_sync2 <= fd_main_tcr_set_time_sync1;
    regs_o.tcr_set_time_o <= fd_main_tcr_set_time_sync2 and (not fd_main_tcr_set_time_sync1);
  end if;
end process;


-- TAI seconds (MSB)
-- asynchronous std_logic_vector register : TAI seconds (MSB) (type RW/WO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_tm_sech_lw_s0 <= '0';
    fd_main_tm_sech_lw_s1 <= '0';
    fd_main_tm_sech_lw_s2 <= '0';
    regs_o.tm_sech_o <= "00000000";
    regs_o.tm_sech_load_o <= '0';
    fd_main_tm_sech_int_read <= "00000000";
  elsif rising_edge(clk_ref_i) then
    fd_main_tm_sech_lw_s0 <= fd_main_tm_sech_lw;
    fd_main_tm_sech_lw_s1 <= fd_main_tm_sech_lw_s0;
    fd_main_tm_sech_lw_s2 <= fd_main_tm_sech_lw_s1;
    if ((fd_main_tm_sech_lw_s2 = '0') and (fd_main_tm_sech_lw_s1 = '1')) then
      if (fd_main_tm_sech_rwsel = '1') then
        regs_o.tm_sech_o <= fd_main_tm_sech_int_write;
        regs_o.tm_sech_load_o <= '1';
      else
        regs_o.tm_sech_load_o <= '0';
        fd_main_tm_sech_int_read <= regs_i.tm_sech_i;
      end if;
    else
      regs_o.tm_sech_load_o <= '0';
    end if;
  end if;
end process;


-- TAI seconds (LSB)
-- asynchronous std_logic_vector register : TAI seconds (LSB) (type RW/WO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_tm_secl_lw_s0 <= '0';
    fd_main_tm_secl_lw_s1 <= '0';
    fd_main_tm_secl_lw_s2 <= '0';
    regs_o.tm_secl_o <= "00000000000000000000000000000000";
    regs_o.tm_secl_load_o <= '0';
    fd_main_tm_secl_int_read <= "00000000000000000000000000000000";
  elsif rising_edge(clk_ref_i) then
    fd_main_tm_secl_lw_s0 <= fd_main_tm_secl_lw;
    fd_main_tm_secl_lw_s1 <= fd_main_tm_secl_lw_s0;
    fd_main_tm_secl_lw_s2 <= fd_main_tm_secl_lw_s1;
    if ((fd_main_tm_secl_lw_s2 = '0') and (fd_main_tm_secl_lw_s1 = '1')) then
      if (fd_main_tm_secl_rwsel = '1') then
        regs_o.tm_secl_o <= fd_main_tm_secl_int_write;
        regs_o.tm_secl_load_o <= '1';
      else
        regs_o.tm_secl_load_o <= '0';
        fd_main_tm_secl_int_read <= regs_i.tm_secl_i;
      end if;
    else
      regs_o.tm_secl_load_o <= '0';
    end if;
  end if;
end process;


-- Reference clock cycles (0...124999999)
-- asynchronous std_logic_vector register : Reference clock cycles (0...124999999) (type RW/WO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_tm_cycles_lw_s0 <= '0';
    fd_main_tm_cycles_lw_s1 <= '0';
    fd_main_tm_cycles_lw_s2 <= '0';
    regs_o.tm_cycles_o <= "0000000000000000000000000000";
    regs_o.tm_cycles_load_o <= '0';
    fd_main_tm_cycles_int_read <= "0000000000000000000000000000";
  elsif rising_edge(clk_ref_i) then
    fd_main_tm_cycles_lw_s0 <= fd_main_tm_cycles_lw;
    fd_main_tm_cycles_lw_s1 <= fd_main_tm_cycles_lw_s0;
    fd_main_tm_cycles_lw_s2 <= fd_main_tm_cycles_lw_s1;
    if ((fd_main_tm_cycles_lw_s2 = '0') and (fd_main_tm_cycles_lw_s1 = '1')) then
      if (fd_main_tm_cycles_rwsel = '1') then
        regs_o.tm_cycles_o <= fd_main_tm_cycles_int_write;
        regs_o.tm_cycles_load_o <= '1';
      else
        regs_o.tm_cycles_load_o <= '0';
        fd_main_tm_cycles_int_read <= regs_i.tm_cycles_i;
      end if;
    else
      regs_o.tm_cycles_load_o <= '0';
    end if;
  end if;
end process;


-- TDC Data
-- asynchronous std_logic_vector register : TDC Data (type RW/WO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_tdr_lw_s0 <= '0';
    fd_main_tdr_lw_s1 <= '0';
    fd_main_tdr_lw_s2 <= '0';
    regs_o.tdr_o <= "0000000000000000000000000000";
    regs_o.tdr_load_o <= '0';
    fd_main_tdr_int_read <= "0000000000000000000000000000";
  elsif rising_edge(clk_ref_i) then
    fd_main_tdr_lw_s0 <= fd_main_tdr_lw;
    fd_main_tdr_lw_s1 <= fd_main_tdr_lw_s0;
    fd_main_tdr_lw_s2 <= fd_main_tdr_lw_s1;
    if ((fd_main_tdr_lw_s2 = '0') and (fd_main_tdr_lw_s1 = '1')) then
      if (fd_main_tdr_rwsel = '1') then
        regs_o.tdr_o <= fd_main_tdr_int_write;
        regs_o.tdr_load_o <= '1';
      else
        regs_o.tdr_load_o <= '0';
        fd_main_tdr_int_read <= regs_i.tdr_i;
      end if;
    else
      regs_o.tdr_load_o <= '0';
    end if;
  end if;
end process;


-- Write to TDC
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.tdcsr_write_o <= '0';
    fd_main_tdcsr_write_sync0 <= '0';
    fd_main_tdcsr_write_sync1 <= '0';
    fd_main_tdcsr_write_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_tdcsr_write_sync0 <= fd_main_tdcsr_write_int;
    fd_main_tdcsr_write_sync1 <= fd_main_tdcsr_write_sync0;
    fd_main_tdcsr_write_sync2 <= fd_main_tdcsr_write_sync1;
    regs_o.tdcsr_write_o <= fd_main_tdcsr_write_sync2 and (not fd_main_tdcsr_write_sync1);
  end if;
end process;


-- Read from TDC
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.tdcsr_read_o <= '0';
    fd_main_tdcsr_read_sync0 <= '0';
    fd_main_tdcsr_read_sync1 <= '0';
    fd_main_tdcsr_read_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_tdcsr_read_sync0 <= fd_main_tdcsr_read_int;
    fd_main_tdcsr_read_sync1 <= fd_main_tdcsr_read_sync0;
    fd_main_tdcsr_read_sync2 <= fd_main_tdcsr_read_sync1;
    regs_o.tdcsr_read_o <= fd_main_tdcsr_read_sync2 and (not fd_main_tdcsr_read_sync1);
  end if;
end process;


-- Empty flag
-- synchronizer chain for field : Empty flag (type RO/WO, clk_ref_i -> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_tdcsr_empty_sync0 <= '0';
    fd_main_tdcsr_empty_sync1 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_tdcsr_empty_sync0 <= regs_i.tdcsr_empty_i;
    fd_main_tdcsr_empty_sync1 <= fd_main_tdcsr_empty_sync0;
  end if;
end process;


-- Stop enable
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.tdcsr_stop_en_o <= '0';
    fd_main_tdcsr_stop_en_sync0 <= '0';
    fd_main_tdcsr_stop_en_sync1 <= '0';
    fd_main_tdcsr_stop_en_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_tdcsr_stop_en_sync0 <= fd_main_tdcsr_stop_en_int;
    fd_main_tdcsr_stop_en_sync1 <= fd_main_tdcsr_stop_en_sync0;
    fd_main_tdcsr_stop_en_sync2 <= fd_main_tdcsr_stop_en_sync1;
    regs_o.tdcsr_stop_en_o <= fd_main_tdcsr_stop_en_sync2 and (not fd_main_tdcsr_stop_en_sync1);
  end if;
end process;


-- Start disable
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.tdcsr_start_dis_o <= '0';
    fd_main_tdcsr_start_dis_sync0 <= '0';
    fd_main_tdcsr_start_dis_sync1 <= '0';
    fd_main_tdcsr_start_dis_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_tdcsr_start_dis_sync0 <= fd_main_tdcsr_start_dis_int;
    fd_main_tdcsr_start_dis_sync1 <= fd_main_tdcsr_start_dis_sync0;
    fd_main_tdcsr_start_dis_sync2 <= fd_main_tdcsr_start_dis_sync1;
    regs_o.tdcsr_start_dis_o <= fd_main_tdcsr_start_dis_sync2 and (not fd_main_tdcsr_start_dis_sync1);
  end if;
end process;


-- Start enable
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.tdcsr_start_en_o <= '0';
    fd_main_tdcsr_start_en_sync0 <= '0';
    fd_main_tdcsr_start_en_sync1 <= '0';
    fd_main_tdcsr_start_en_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_tdcsr_start_en_sync0 <= fd_main_tdcsr_start_en_int;
    fd_main_tdcsr_start_en_sync1 <= fd_main_tdcsr_start_en_sync0;
    fd_main_tdcsr_start_en_sync2 <= fd_main_tdcsr_start_en_sync1;
    regs_o.tdcsr_start_en_o <= fd_main_tdcsr_start_en_sync2 and (not fd_main_tdcsr_start_en_sync1);
  end if;
end process;


-- Stop disable
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.tdcsr_stop_dis_o <= '0';
    fd_main_tdcsr_stop_dis_sync0 <= '0';
    fd_main_tdcsr_stop_dis_sync1 <= '0';
    fd_main_tdcsr_stop_dis_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_tdcsr_stop_dis_sync0 <= fd_main_tdcsr_stop_dis_int;
    fd_main_tdcsr_stop_dis_sync1 <= fd_main_tdcsr_stop_dis_sync0;
    fd_main_tdcsr_stop_dis_sync2 <= fd_main_tdcsr_stop_dis_sync1;
    regs_o.tdcsr_stop_dis_o <= fd_main_tdcsr_stop_dis_sync2 and (not fd_main_tdcsr_stop_dis_sync1);
  end if;
end process;


-- Pulse <code>Alutrigger</code> line
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.tdcsr_alutrig_o <= '0';
    fd_main_tdcsr_alutrig_sync0 <= '0';
    fd_main_tdcsr_alutrig_sync1 <= '0';
    fd_main_tdcsr_alutrig_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_tdcsr_alutrig_sync0 <= fd_main_tdcsr_alutrig_int;
    fd_main_tdcsr_alutrig_sync1 <= fd_main_tdcsr_alutrig_sync0;
    fd_main_tdcsr_alutrig_sync2 <= fd_main_tdcsr_alutrig_sync1;
    regs_o.tdcsr_alutrig_o <= fd_main_tdcsr_alutrig_sync2 and (not fd_main_tdcsr_alutrig_sync1);
  end if;
end process;


-- IDELAY CE (pulse)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.tdcsr_idelay_ce_o <= '0';
    fd_main_tdcsr_idelay_ce_sync0 <= '0';
    fd_main_tdcsr_idelay_ce_sync1 <= '0';
    fd_main_tdcsr_idelay_ce_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_tdcsr_idelay_ce_sync0 <= fd_main_tdcsr_idelay_ce_int;
    fd_main_tdcsr_idelay_ce_sync1 <= fd_main_tdcsr_idelay_ce_sync0;
    fd_main_tdcsr_idelay_ce_sync2 <= fd_main_tdcsr_idelay_ce_sync1;
    regs_o.tdcsr_idelay_ce_o <= fd_main_tdcsr_idelay_ce_sync2 and (not fd_main_tdcsr_idelay_ce_sync1);
  end if;
end process;


-- Generate calibration pulses (type 1 calibration)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.calr_cal_pulse_o <= '0';
    fd_main_calr_cal_pulse_sync0 <= '0';
    fd_main_calr_cal_pulse_sync1 <= '0';
    fd_main_calr_cal_pulse_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_calr_cal_pulse_sync0 <= fd_main_calr_cal_pulse_int;
    fd_main_calr_cal_pulse_sync1 <= fd_main_calr_cal_pulse_sync0;
    fd_main_calr_cal_pulse_sync2 <= fd_main_calr_cal_pulse_sync1;
    regs_o.calr_cal_pulse_o <= fd_main_calr_cal_pulse_sync2 and (not fd_main_calr_cal_pulse_sync1);
  end if;
end process;


-- PPS calibration output enable.
-- synchronizer chain for field : PPS calibration output enable. (type RW/RO, clk_sys_i <-> clk_ref_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.calr_cal_pps_o <= '0';
    fd_main_calr_cal_pps_sync0 <= '0';
    fd_main_calr_cal_pps_sync1 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_calr_cal_pps_sync0 <= fd_main_calr_cal_pps_int;
    fd_main_calr_cal_pps_sync1 <= fd_main_calr_cal_pps_sync0;
    regs_o.calr_cal_pps_o <= fd_main_calr_cal_pps_sync1;
  end if;
end process;


-- Produce DDMTD calibration pattern (type 2 calibration)
regs_o.calr_cal_dmtd_o <= fd_main_calr_cal_dmtd_int;
-- Calibration pulse output select/mask
-- asynchronous std_logic_vector register : Calibration pulse output select/mask (type RW/RO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_calr_psel_swb_s0 <= '0';
    fd_main_calr_psel_swb_s1 <= '0';
    fd_main_calr_psel_swb_s2 <= '0';
    regs_o.calr_psel_o <= "0000";
  elsif rising_edge(clk_ref_i) then
    fd_main_calr_psel_swb_s0 <= fd_main_calr_psel_swb;
    fd_main_calr_psel_swb_s1 <= fd_main_calr_psel_swb_s0;
    fd_main_calr_psel_swb_s2 <= fd_main_calr_psel_swb_s1;
    if ((fd_main_calr_psel_swb_s2 = '0') and (fd_main_calr_psel_swb_s1 = '1')) then
      regs_o.calr_psel_o <= fd_main_calr_psel_int;
    end if;
  end if;
end process;


-- DMTD Tag
-- DMTD Tag Ready
-- DMTD Tag
-- DMTD Tag Ready
-- ADSFR Value
-- asynchronous std_logic_vector register : ADSFR Value (type RW/RO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_adsfr_swb_s0 <= '0';
    fd_main_adsfr_swb_s1 <= '0';
    fd_main_adsfr_swb_s2 <= '0';
    regs_o.adsfr_o <= "000000000000000000";
  elsif rising_edge(clk_ref_i) then
    fd_main_adsfr_swb_s0 <= fd_main_adsfr_swb;
    fd_main_adsfr_swb_s1 <= fd_main_adsfr_swb_s0;
    fd_main_adsfr_swb_s2 <= fd_main_adsfr_swb_s1;
    if ((fd_main_adsfr_swb_s2 = '0') and (fd_main_adsfr_swb_s1 = '1')) then
      regs_o.adsfr_o <= fd_main_adsfr_int;
    end if;
  end if;
end process;


-- Coarse threshold
-- asynchronous std_logic_vector register : Coarse threshold (type RW/RO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_atmcr_c_thr_swb_s0 <= '0';
    fd_main_atmcr_c_thr_swb_s1 <= '0';
    fd_main_atmcr_c_thr_swb_s2 <= '0';
    regs_o.atmcr_c_thr_o <= "00000000";
  elsif rising_edge(clk_ref_i) then
    fd_main_atmcr_c_thr_swb_s0 <= fd_main_atmcr_c_thr_swb;
    fd_main_atmcr_c_thr_swb_s1 <= fd_main_atmcr_c_thr_swb_s0;
    fd_main_atmcr_c_thr_swb_s2 <= fd_main_atmcr_c_thr_swb_s1;
    if ((fd_main_atmcr_c_thr_swb_s2 = '0') and (fd_main_atmcr_c_thr_swb_s1 = '1')) then
      regs_o.atmcr_c_thr_o <= fd_main_atmcr_c_thr_int;
    end if;
  end if;
end process;


-- Fine threshold
-- asynchronous std_logic_vector register : Fine threshold (type RW/RO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_atmcr_f_thr_swb_s0 <= '0';
    fd_main_atmcr_f_thr_swb_s1 <= '0';
    fd_main_atmcr_f_thr_swb_s2 <= '0';
    regs_o.atmcr_f_thr_o <= "00000000000000000000000";
  elsif rising_edge(clk_ref_i) then
    fd_main_atmcr_f_thr_swb_s0 <= fd_main_atmcr_f_thr_swb;
    fd_main_atmcr_f_thr_swb_s1 <= fd_main_atmcr_f_thr_swb_s0;
    fd_main_atmcr_f_thr_swb_s2 <= fd_main_atmcr_f_thr_swb_s1;
    if ((fd_main_atmcr_f_thr_swb_s2 = '0') and (fd_main_atmcr_f_thr_swb_s1 = '1')) then
      regs_o.atmcr_f_thr_o <= fd_main_atmcr_f_thr_int;
    end if;
  end if;
end process;


-- Start Offset
-- asynchronous std_logic_vector register : Start Offset (type RW/RO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_asor_offset_swb_s0 <= '0';
    fd_main_asor_offset_swb_s1 <= '0';
    fd_main_asor_offset_swb_s2 <= '0';
    regs_o.asor_offset_o <= "00000000000000000000000";
  elsif rising_edge(clk_ref_i) then
    fd_main_asor_offset_swb_s0 <= fd_main_asor_offset_swb;
    fd_main_asor_offset_swb_s1 <= fd_main_asor_offset_swb_s0;
    fd_main_asor_offset_swb_s2 <= fd_main_asor_offset_swb_s1;
    if ((fd_main_asor_offset_swb_s2 = '0') and (fd_main_asor_offset_swb_s1 = '1')) then
      regs_o.asor_offset_o <= fd_main_asor_offset_int;
    end if;
  end if;
end process;


-- Number of raw events.
-- asynchronous std_logic_vector register : Number of raw events. (type RO/WO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_iecraw_lwb_s0 <= '0';
    fd_main_iecraw_lwb_s1 <= '0';
    fd_main_iecraw_lwb_s2 <= '0';
    fd_main_iecraw_int <= "00000000000000000000000000000000";
  elsif rising_edge(clk_ref_i) then
    fd_main_iecraw_lwb_s0 <= fd_main_iecraw_lwb;
    fd_main_iecraw_lwb_s1 <= fd_main_iecraw_lwb_s0;
    fd_main_iecraw_lwb_s2 <= fd_main_iecraw_lwb_s1;
    if ((fd_main_iecraw_lwb_s1 = '1') and (fd_main_iecraw_lwb_s2 = '0')) then
      fd_main_iecraw_int <= regs_i.iecraw_i;
    end if;
  end if;
end process;


-- Number of tagged events
-- asynchronous std_logic_vector register : Number of tagged events (type RO/WO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_iectag_lwb_s0 <= '0';
    fd_main_iectag_lwb_s1 <= '0';
    fd_main_iectag_lwb_s2 <= '0';
    fd_main_iectag_int <= "00000000000000000000000000000000";
  elsif rising_edge(clk_ref_i) then
    fd_main_iectag_lwb_s0 <= fd_main_iectag_lwb;
    fd_main_iectag_lwb_s1 <= fd_main_iectag_lwb_s0;
    fd_main_iectag_lwb_s2 <= fd_main_iectag_lwb_s1;
    if ((fd_main_iectag_lwb_s1 = '1') and (fd_main_iectag_lwb_s2 = '0')) then
      fd_main_iectag_int <= regs_i.iectag_i;
    end if;
  end if;
end process;


-- Reset stats
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.iepd_rst_stat_o <= '0';
    fd_main_iepd_rst_stat_sync0 <= '0';
    fd_main_iepd_rst_stat_sync1 <= '0';
    fd_main_iepd_rst_stat_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_iepd_rst_stat_sync0 <= fd_main_iepd_rst_stat_int;
    fd_main_iepd_rst_stat_sync1 <= fd_main_iepd_rst_stat_sync0;
    fd_main_iepd_rst_stat_sync2 <= fd_main_iepd_rst_stat_sync1;
    regs_o.iepd_rst_stat_o <= fd_main_iepd_rst_stat_sync2 and (not fd_main_iepd_rst_stat_sync1);
  end if;
end process;


-- Processing delay
-- asynchronous std_logic_vector register : Processing delay (type RO/WO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_iepd_pdelay_lwb_s0 <= '0';
    fd_main_iepd_pdelay_lwb_s1 <= '0';
    fd_main_iepd_pdelay_lwb_s2 <= '0';
    fd_main_iepd_pdelay_int <= "00000000";
  elsif rising_edge(clk_ref_i) then
    fd_main_iepd_pdelay_lwb_s0 <= fd_main_iepd_pdelay_lwb;
    fd_main_iepd_pdelay_lwb_s1 <= fd_main_iepd_pdelay_lwb_s0;
    fd_main_iepd_pdelay_lwb_s2 <= fd_main_iepd_pdelay_lwb_s1;
    if ((fd_main_iepd_pdelay_lwb_s1 = '1') and (fd_main_iepd_pdelay_lwb_s2 = '0')) then
      fd_main_iepd_pdelay_int <= regs_i.iepd_pdelay_i;
    end if;
  end if;
end process;


-- Data
regs_o.scr_data_o <= wrdata_reg(23 downto 0);
-- Select DAC
regs_o.scr_sel_dac_o <= fd_main_scr_sel_dac_int;
-- Select PLL
regs_o.scr_sel_pll_o <= fd_main_scr_sel_pll_int;
-- Select GPIO
regs_o.scr_sel_gpio_o <= fd_main_scr_sel_gpio_int;
-- Ready flag
-- Clock Polarity
regs_o.scr_cpol_o <= fd_main_scr_cpol_int;
-- Transfer Start
process (clk_sys_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_scr_start_dly0 <= '0';
    regs_o.scr_start_o <= '0';
  elsif rising_edge(clk_sys_i) then
    fd_main_scr_start_dly0 <= fd_main_scr_start_int;
    regs_o.scr_start_o <= fd_main_scr_start_int and (not fd_main_scr_start_dly0);
  end if;
end process;


-- Frequency
-- asynchronous std_logic_vector register : Frequency (type RO/WO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_rcrr_lwb_s0 <= '0';
    fd_main_rcrr_lwb_s1 <= '0';
    fd_main_rcrr_lwb_s2 <= '0';
    fd_main_rcrr_int <= "00000000000000000000000000000000";
  elsif rising_edge(clk_ref_i) then
    fd_main_rcrr_lwb_s0 <= fd_main_rcrr_lwb;
    fd_main_rcrr_lwb_s1 <= fd_main_rcrr_lwb_s0;
    fd_main_rcrr_lwb_s2 <= fd_main_rcrr_lwb_s1;
    if ((fd_main_rcrr_lwb_s1 = '1') and (fd_main_rcrr_lwb_s2 = '0')) then
      fd_main_rcrr_int <= regs_i.rcrr_i;
    end if;
  end if;
end process;


-- Channel mask
-- asynchronous std_logic_vector register : Channel mask (type RW/RO, clk_ref_i <-> clk_sys_i)
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_tsbcr_chan_mask_swb_s0 <= '0';
    fd_main_tsbcr_chan_mask_swb_s1 <= '0';
    fd_main_tsbcr_chan_mask_swb_s2 <= '0';
    regs_o.tsbcr_chan_mask_o <= "00000";
  elsif rising_edge(clk_ref_i) then
    fd_main_tsbcr_chan_mask_swb_s0 <= fd_main_tsbcr_chan_mask_swb;
    fd_main_tsbcr_chan_mask_swb_s1 <= fd_main_tsbcr_chan_mask_swb_s0;
    fd_main_tsbcr_chan_mask_swb_s2 <= fd_main_tsbcr_chan_mask_swb_s1;
    if ((fd_main_tsbcr_chan_mask_swb_s2 = '0') and (fd_main_tsbcr_chan_mask_swb_s1 = '1')) then
      regs_o.tsbcr_chan_mask_o <= fd_main_tsbcr_chan_mask_int;
    end if;
  end if;
end process;


-- Buffer enable
regs_o.tsbcr_enable_o <= fd_main_tsbcr_enable_int;
-- Buffer purge
process (clk_sys_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_tsbcr_purge_dly0 <= '0';
    regs_o.tsbcr_purge_o <= '0';
  elsif rising_edge(clk_sys_i) then
    fd_main_tsbcr_purge_dly0 <= fd_main_tsbcr_purge_int;
    regs_o.tsbcr_purge_o <= fd_main_tsbcr_purge_int and (not fd_main_tsbcr_purge_dly0);
  end if;
end process;


-- Reset timestamp sequence number
process (clk_ref_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    regs_o.tsbcr_rst_seq_o <= '0';
    fd_main_tsbcr_rst_seq_sync0 <= '0';
    fd_main_tsbcr_rst_seq_sync1 <= '0';
    fd_main_tsbcr_rst_seq_sync2 <= '0';
  elsif rising_edge(clk_ref_i) then
    fd_main_tsbcr_rst_seq_sync0 <= fd_main_tsbcr_rst_seq_int;
    fd_main_tsbcr_rst_seq_sync1 <= fd_main_tsbcr_rst_seq_sync0;
    fd_main_tsbcr_rst_seq_sync2 <= fd_main_tsbcr_rst_seq_sync1;
    regs_o.tsbcr_rst_seq_o <= fd_main_tsbcr_rst_seq_sync2 and (not fd_main_tsbcr_rst_seq_sync1);
  end if;
end process;


-- Buffer full
-- Buffer empty
-- Buffer entries count
-- RAW readout mode enable
regs_o.tsbcr_raw_o <= fd_main_tsbcr_raw_int;
-- IRQ timeout [milliseconds]
regs_o.tsbir_timeout_o <= fd_main_tsbir_timeout_int;
-- Interrupt threshold
regs_o.tsbir_threshold_o <= fd_main_tsbir_threshold_int;
-- Timestamps TAI Seconds (bits 39-32)
-- Timestamps TAI Seconds (bits 31-0)
-- Timestamps cycles count (in 8 ns ticks)
-- Channel ID
-- Fine Value (in phase units)
-- Timestamp Sequence ID
-- SCL Line out
regs_o.i2cr_scl_out_o <= fd_main_i2cr_scl_out_int;
-- SDA Line out
regs_o.i2cr_sda_out_o <= fd_main_i2cr_sda_out_int;
-- SCL Line in
-- SDA Line in
-- VCXO Frequency
-- Peltier PWM drive
regs_o.tder2_pelt_drive_o <= fd_main_tder2_pelt_drive_int;
-- Debug value
-- Advance buffer readout
process (clk_sys_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    fd_main_tsbr_advance_adv_dly0 <= '0';
    regs_o.tsbr_advance_adv_o <= '0';
  elsif rising_edge(clk_sys_i) then
    fd_main_tsbr_advance_adv_dly0 <= fd_main_tsbr_advance_adv_int;
    regs_o.tsbr_advance_adv_o <= fd_main_tsbr_advance_adv_int and (not fd_main_tsbr_advance_adv_dly0);
  end if;
end process;


-- Slot ID
-- Number of delay line taps.
regs_o.iodelay_adj_n_taps_o <= wrdata_reg(7 downto 0);
-- extra code for reg/fifo/mem: Interrupt disable register
eic_idr_int(2 downto 0) <= wrdata_reg(2 downto 0);
-- extra code for reg/fifo/mem: Interrupt enable register
eic_ier_int(2 downto 0) <= wrdata_reg(2 downto 0);
-- extra code for reg/fifo/mem: Interrupt status register
eic_isr_clear_int(2 downto 0) <= wrdata_reg(2 downto 0);
-- extra code for reg/fifo/mem: IRQ_CONTROLLER
eic_irq_controller_inst : wbgen2_eic
  generic map (
    g_num_interrupts     => 3,
    g_irq00_mode         => 3,
    g_irq01_mode         => 0,
    g_irq02_mode         => 0,
    g_irq03_mode         => 0,
    g_irq04_mode         => 0,
    g_irq05_mode         => 0,
    g_irq06_mode         => 0,
    g_irq07_mode         => 0,
    g_irq08_mode         => 0,
    g_irq09_mode         => 0,
    g_irq0a_mode         => 0,
    g_irq0b_mode         => 0,
    g_irq0c_mode         => 0,
    g_irq0d_mode         => 0,
    g_irq0e_mode         => 0,
    g_irq0f_mode         => 0,
    g_irq10_mode         => 0,
    g_irq11_mode         => 0,
    g_irq12_mode         => 0,
    g_irq13_mode         => 0,
    g_irq14_mode         => 0,
    g_irq15_mode         => 0,
    g_irq16_mode         => 0,
    g_irq17_mode         => 0,
    g_irq18_mode         => 0,
    g_irq19_mode         => 0,
    g_irq1a_mode         => 0,
    g_irq1b_mode         => 0,
    g_irq1c_mode         => 0,
    g_irq1d_mode         => 0,
    g_irq1e_mode         => 0,
    g_irq1f_mode         => 0
  )
  port map (
    clk_i                => clk_sys_i,
    rst_n_i              => rst_n_i,
    irq_i                => irq_inputs_vector_int,
    irq_ack_o            => eic_irq_ack_int,
    reg_imr_o            => eic_imr_int,
    reg_ier_i            => eic_ier_int,
    reg_ier_wr_stb_i     => eic_ier_write_int,
    reg_idr_i            => eic_idr_int,
    reg_idr_wr_stb_i     => eic_idr_write_int,
    reg_isr_o            => eic_isr_status_int,
    reg_isr_i            => eic_isr_clear_int,
    reg_isr_wr_stb_i     => eic_isr_write_int,
    wb_irq_o             => wb_int_o
  );

irq_inputs_vector_int(0) <= irq_ts_buf_notempty_i;
irq_inputs_vector_int(1) <= irq_dmtd_spll_i;
irq_inputs_vector_int(2) <= irq_sync_status_i;
rwaddr_reg <= wb_adr_i;
wb_stall_o <= (not ack_sreg(0)) and (wb_stb_i and wb_cyc_i);
wb_err_o <= '0';
wb_rty_o <= '0';
-- ACK signal generation. Just pass the LSB of ACK counter.
wb_ack_o <= ack_sreg(0);
end syn;
